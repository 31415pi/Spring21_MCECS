Char
Code
Hex Binary a b c d e f g

Special Characters
Char
Code
Hex Binary a b c d e f g Description
function logic [7:0] BtS ( input logic [4:0] binaryvalues ) ;


0 00 00000 1 1 1 1 1 1 0
1 01 00001 0 0 0 0 1 1 0
2 02 00010 1 1 0 1 1 0 1
3 03 00011 1 1 1 1 0 0 1
4 04 00100 0 1 1 0 0 1 1
5 05 00101 1 0 1 1 0 1 1
6 06 00110 1 0 1 1 1 1 1
7 07 00111 1 1 1 0 0 0 0
8 08 01000 1 1 1 1 1 1 1
9 09 01001 1 1 1 1 0 1 1
10 0A 01010 1 1 1 0 1 1 1
11 0B 01011 0 0 1 1 1 1 1
12 0C 01100 1 0 0 1 1 1 0
13 0D 01101 0 1 1 1 1 0 1
14 0E 01110 1 0 0 1 1 1 1
15 0F 01111 1 0 0 0 1 1 1
16 10 10000 1 0 0 0 0 0 0 Segment a
17 11 00001 0 1 0 0 0 0 0 Segment b
18 12 10010 0 0 1 0 0 0 0 Segment c
19 13 10011 0 0 0 1 0 0 0 Segment d
20 14 10100 0 0 0 0 1 0 0 Segment e
21 15 10101 0 0 0 0 0 1 0 Segment f
22 16 10110 0 0 0 0 0 0 1 Segment g
23 17 10111 0 0 0 0 0 0 0 BLANK
24 18 11000 0 1 1 0 1 1 1 Upper case H
25 19 11001 0 0 0 1 1 1 0 Upper case L
26 1A 11010 1 1 1 0 1 1 1 Upper case R
27 1B 11011 0 0 0 0 1 1 0 Lower case L
28 1C 11100 0 0 0 0 1 0 1 Lower case R
29 1D 11101 0 0 0 0 0 0 0 BLANK
30 1E 11110 0 0 0 0 0 0 0 BLANK
31 1F 11111 0 0 0 0 0 0 0 BLANK